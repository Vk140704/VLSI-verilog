module not_gate (
    input a,   // Input A
    output y   // Output Y
);
    assign y = ~a;  // NOT operation
endmodule

